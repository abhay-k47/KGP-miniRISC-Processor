`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:28:26 11/09/2022 
// Design Name: 
// Module Name:    Decoder 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Decoder(
    input [31:0] in,
    output reg [31:0] out
    );
	always@(*)begin
		case(in)
			32'b00000000000000000000000000000001: out <= {{27{1'b0}},5'd0};
			32'b00000000000000000000000000000010: out <= {{27{1'b0}},5'd1};
			32'b00000000000000000000000000000100: out <= {{27{1'b0}},5'd2};
			32'b00000000000000000000000000001000: out <= {{27{1'b0}},5'd3};
			32'b00000000000000000000000000010000: out <= {{27{1'b0}},5'd4};
			32'b00000000000000000000000000100000: out <= {{27{1'b0}},5'd5};
			32'b00000000000000000000000001000000: out <= {{27{1'b0}},5'd6};
			32'b00000000000000000000000010000000: out <= {{27{1'b0}},5'd7};
			32'b00000000000000000000000100000000: out <= {{27{1'b0}},5'd8};
			32'b00000000000000000000001000000000: out <= {{27{1'b0}},5'd9};
			32'b00000000000000000000010000000000: out <= {{27{1'b0}},5'd10};
			32'b00000000000000000000100000000000: out <= {{27{1'b0}},5'd11};
			32'b00000000000000000001000000000000: out <= {{27{1'b0}},5'd12};
			32'b00000000000000000010000000000000: out <= {{27{1'b0}},5'd13};
			32'b00000000000000000100000000000000: out <= {{27{1'b0}},5'd14};
			32'b00000000000000001000000000000000: out <= {{27{1'b0}},5'd15};
			32'b00000000000000010000000000000000: out <= {{27{1'b0}},5'd16};
			32'b00000000000000100000000000000000: out <= {{27{1'b0}},5'd17};
			32'b00000000000001000000000000000000: out <= {{27{1'b0}},5'd18};
			32'b00000000000010000000000000000000: out <= {{27{1'b0}},5'd19};
			32'b00000000000100000000000000000000: out <= {{27{1'b0}},5'd20};
			32'b00000000001000000000000000000000: out <= {{27{1'b0}},5'd21};
			32'b00000000010000000000000000000000: out <= {{27{1'b0}},5'd22};
			32'b00000000100000000000000000000000: out <= {{27{1'b0}},5'd23};
			32'b00000001000000000000000000000000: out <= {{27{1'b0}},5'd24};
			32'b00000010000000000000000000000000: out <= {{27{1'b0}},5'd25};
			32'b00000100000000000000000000000000: out <= {{27{1'b0}},5'd26};
			32'b00001000000000000000000000000000: out <= {{27{1'b0}},5'd27};
			32'b00010000000000000000000000000000: out <= {{27{1'b0}},5'd28};
			32'b00100000000000000000000000000000: out <= {{27{1'b0}},5'd29};
			32'b01000000000000000000000000000000: out <= {{27{1'b0}},5'd30};
			32'b10000000000000000000000000000000: out <= {{27{1'b0}},5'd31};
			default: out <= {32{1'b1}};
		endcase
	end

endmodule
